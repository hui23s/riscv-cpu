`include "../chip_param.v"

module core_ifu (
    input wire clk_i,
    input wire rst_n_i
  );

  // do nothing here!

endmodule
